//
//
//
module i2c_extender (
input sda,
input scl,
output scl,
output sda1,
output sda2,
);

endmodule
